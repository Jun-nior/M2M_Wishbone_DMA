package DMA_CSR_rtl_pkg;
  localparam int SOURCE_ADDR_REG_BYTE_WIDTH = 4;
  localparam int SOURCE_ADDR_REG_BYTE_SIZE = 4;
  localparam bit [4:0] SOURCE_ADDR_REG_BYTE_OFFSET = 5'h00;
  localparam int SOURCE_ADDR_REG_ADDR_BIT_WIDTH = 32;
  localparam bit [31:0] SOURCE_ADDR_REG_ADDR_BIT_MASK = 32'hffffffff;
  localparam int SOURCE_ADDR_REG_ADDR_BIT_OFFSET = 0;
  localparam int DEST_ADDR_REG_BYTE_WIDTH = 4;
  localparam int DEST_ADDR_REG_BYTE_SIZE = 4;
  localparam bit [4:0] DEST_ADDR_REG_BYTE_OFFSET = 5'h04;
  localparam int DEST_ADDR_REG_ADDR_BIT_WIDTH = 32;
  localparam bit [31:0] DEST_ADDR_REG_ADDR_BIT_MASK = 32'hffffffff;
  localparam int DEST_ADDR_REG_ADDR_BIT_OFFSET = 0;
  localparam int LENGTH_REG_BYTE_WIDTH = 4;
  localparam int LENGTH_REG_BYTE_SIZE = 4;
  localparam bit [4:0] LENGTH_REG_BYTE_OFFSET = 5'h08;
  localparam int LENGTH_REG_LEN_BIT_WIDTH = 16;
  localparam bit [15:0] LENGTH_REG_LEN_BIT_MASK = 16'hffff;
  localparam int LENGTH_REG_LEN_BIT_OFFSET = 0;
  localparam int CONTROL_REG_BYTE_WIDTH = 4;
  localparam int CONTROL_REG_BYTE_SIZE = 4;
  localparam bit [4:0] CONTROL_REG_BYTE_OFFSET = 5'h0c;
  localparam int CONTROL_REG_GO_BIT_WIDTH = 1;
  localparam bit CONTROL_REG_GO_BIT_MASK = 1'h1;
  localparam int CONTROL_REG_GO_BIT_OFFSET = 0;
  localparam int CONTROL_REG_IE_BIT_WIDTH = 1;
  localparam bit CONTROL_REG_IE_BIT_MASK = 1'h1;
  localparam int CONTROL_REG_IE_BIT_OFFSET = 1;
  localparam int STATUS_REG_BYTE_WIDTH = 4;
  localparam int STATUS_REG_BYTE_SIZE = 4;
  localparam bit [4:0] STATUS_REG_BYTE_OFFSET = 5'h10;
  localparam int STATUS_REG_BUSY_BIT_WIDTH = 1;
  localparam bit STATUS_REG_BUSY_BIT_MASK = 1'h1;
  localparam int STATUS_REG_BUSY_BIT_OFFSET = 0;
  localparam int STATUS_REG_DONE_IF_BIT_WIDTH = 1;
  localparam bit STATUS_REG_DONE_IF_BIT_MASK = 1'h1;
  localparam int STATUS_REG_DONE_IF_BIT_OFFSET = 16;
endpackage
